module seg7(output reg [6:0]s,input [3:]b);
 always @ (b)
 begin
 s=7'b0000000;
 b=4'b0000;
 case(b)
 4'b0000:s=7'b1111110;
 4'b0001:s=7'b0110000;
 4'b0010:s=7'b1101101;
 4'b0000:s=7'b1111110;
 4'b0000:s=7'b1111110;
 4'b0000:s=7'b1111110;
 4'b0000:s=7'b1111110;
 4'b0000:s=7'b1111110;
 4'b0000:s=7'b1111110;
 4'b0000:s=7'b1111110;
 

 
