module sumbytwo(output y,input x2,x1,x0);
	assign y = ~x2;
endmodule
