module four_bit_cla(output cout,[3:0]s,input cin ,[3:0]a,b);
	wire c0,c1,c2;
	wire p0,p1,p2,p3;
	wire g0,g1,g2,g3;
	assign p0=a[0]^b[0];
	assign p1=a[1]^b[1];
	assign p2=a[2]^b[2];
	assign p3=a[3]^b[3];
	assign g0=a[0]&b[0];
	assign g1=a[1]&b[1];
	assign g2=a[2]&b[2];
	assign g3=a[3]&b[3];
	assign c0=(p0&cin)|g0;
	assign c1=(p0&p1&cin)|(p1&g0)|g1;
	assign c2=(p0&p1&p2&cin)|(p1&p2&g0)|(p2&g1)|g2;
	assign cout=(p0&p1&p2&p3&cin)|(p1&p2&p3&g0)|(p2&p3&g1)|(p3&g2)|g3;
	assign s[0]=p0^cin;
	assign s[1]=p1^c0;
	assign s[2]=p2^c1;
	assign s[3]=p3^c2;
endmodule 