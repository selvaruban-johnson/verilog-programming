module orgate(output out, input a, b);
	assign out= a|b;
endmodule 